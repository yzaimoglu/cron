module main

fn main() {
	println('Cron library')
}
